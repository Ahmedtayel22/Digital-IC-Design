module edge_bit_counter (enable, Prescale, CLK, RST, bit_cnt, edge_cnt);
input        enable;
input [5:0]  Prescale;
input        CLK;
input        RST;
output [3:0] bit_cnt;
output [5:0] edge_cnt;

reg [3:0] bit_cnt;
reg [5:0] edge_cnt;

always @(posedge CLK or negedge RST) 
begin
    if(!RST)
    begin
        bit_cnt  <= 4'b0;
        edge_cnt <= 6'b0;
    end
    else if (enable)
    begin
        if (edge_cnt == (Prescale-1)) 
        begin
            bit_cnt <= bit_cnt + 1; 
            edge_cnt <= 0; 
        end
        else edge_cnt <= edge_cnt + 1 ;
    end
    else
    begin
        bit_cnt  <= 4'b0;
        edge_cnt <= 6'b0;
    end
end
endmodule
